library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4067	)	,
(	4063	)	,
(	4059	)	,
(	4055	)	,
(	4052	)	,
(	4048	)	,
(	4044	)	,
(	4040	)	,
(	4036	)	,
(	4032	)	,
(	4029	)	,
(	4025	)	,
(	4021	)	,
(	4017	)	,
(	4013	)	,
(	4010	)	,
(	4006	)	,
(	4002	)	,
(	3998	)	,
(	3994	)	,
(	3991	)	,
(	3987	)	,
(	3983	)	,
(	3979	)	,
(	3975	)	,
(	3972	)	,
(	3968	)	,
(	3964	)	,
(	3960	)	,
(	3957	)	,
(	3953	)	,
(	3949	)	,
(	3945	)	,
(	3941	)	,
(	3938	)	,
(	3934	)	,
(	3930	)	,
(	3926	)	,
(	3923	)	,
(	3919	)	,
(	3915	)	,
(	3911	)	,
(	3908	)	,
(	3904	)	,
(	3900	)	,
(	3897	)	,
(	3893	)	,
(	3889	)	,
(	3885	)	,
(	3882	)	,
(	3878	)	,
(	3874	)	,
(	3870	)	,
(	3867	)	,
(	3863	)	,
(	3859	)	,
(	3856	)	,
(	3852	)	,
(	3848	)	,
(	3845	)	,
(	3841	)	,
(	3837	)	,
(	3833	)	,
(	3830	)	,
(	3826	)	,
(	3822	)	,
(	3819	)	,
(	3815	)	,
(	3811	)	,
(	3808	)	,
(	3804	)	,
(	3800	)	,
(	3797	)	,
(	3793	)	,
(	3789	)	,
(	3786	)	,
(	3782	)	,
(	3778	)	,
(	3775	)	,
(	3771	)	,
(	3768	)	,
(	3764	)	,
(	3760	)	,
(	3757	)	,
(	3753	)	,
(	3749	)	,
(	3746	)	,
(	3742	)	,
(	3738	)	,
(	3735	)	,
(	3731	)	,
(	3728	)	,
(	3724	)	,
(	3720	)	,
(	3717	)	,
(	3713	)	,
(	3710	)	,
(	3706	)	,
(	3702	)	,
(	3699	)	,
(	3695	)	,
(	3692	)	,
(	3688	)	,
(	3684	)	,
(	3681	)	,
(	3677	)	,
(	3674	)	,
(	3670	)	,
(	3667	)	,
(	3663	)	,
(	3659	)	,
(	3656	)	,
(	3652	)	,
(	3649	)	,
(	3645	)	,
(	3642	)	,
(	3638	)	,
(	3634	)	,
(	3631	)	,
(	3627	)	,
(	3624	)	,
(	3620	)	,
(	3617	)	,
(	3613	)	,
(	3610	)	,
(	3606	)	,
(	3603	)	,
(	3599	)	,
(	3596	)	,
(	3592	)	,
(	3589	)	,
(	3585	)	,
(	3582	)	,
(	3578	)	,
(	3575	)	,
(	3571	)	,
(	3567	)	,
(	3564	)	,
(	3560	)	,
(	3557	)	,
(	3554	)	,
(	3550	)	,
(	3547	)	,
(	3543	)	,
(	3540	)	,
(	3536	)	,
(	3533	)	,
(	3529	)	,
(	3526	)	,
(	3522	)	,
(	3519	)	,
(	3515	)	,
(	3512	)	,
(	3508	)	,
(	3505	)	,
(	3501	)	,
(	3498	)	,
(	3494	)	,
(	3491	)	,
(	3488	)	,
(	3484	)	,
(	3481	)	,
(	3477	)	,
(	3474	)	,
(	3470	)	,
(	3467	)	,
(	3464	)	,
(	3460	)	,
(	3457	)	,
(	3453	)	,
(	3450	)	,
(	3446	)	,
(	3443	)	,
(	3440	)	,
(	3436	)	,
(	3433	)	,
(	3429	)	,
(	3426	)	,
(	3423	)	,
(	3419	)	,
(	3416	)	,
(	3412	)	,
(	3409	)	,
(	3406	)	,
(	3402	)	,
(	3399	)	,
(	3395	)	,
(	3392	)	,
(	3389	)	,
(	3385	)	,
(	3382	)	,
(	3379	)	,
(	3375	)	,
(	3372	)	,
(	3368	)	,
(	3365	)	,
(	3362	)	,
(	3358	)	,
(	3355	)	,
(	3352	)	,
(	3348	)	,
(	3345	)	,
(	3342	)	,
(	3338	)	,
(	3335	)	,
(	3332	)	,
(	3328	)	,
(	3325	)	,
(	3322	)	,
(	3318	)	,
(	3315	)	,
(	3312	)	,
(	3308	)	,
(	3305	)	,
(	3302	)	,
(	3298	)	,
(	3295	)	,
(	3292	)	,
(	3288	)	,
(	3285	)	,
(	3282	)	,
(	3279	)	,
(	3275	)	,
(	3272	)	,
(	3269	)	,
(	3265	)	,
(	3262	)	,
(	3259	)	,
(	3256	)	,
(	3252	)	,
(	3249	)	,
(	3246	)	,
(	3242	)	,
(	3239	)	,
(	3236	)	,
(	3233	)	,
(	3229	)	,
(	3226	)	,
(	3223	)	,
(	3220	)	,
(	3216	)	,
(	3213	)	,
(	3210	)	,
(	3207	)	,
(	3203	)	,
(	3200	)	,
(	3197	)	,
(	3194	)	,
(	3190	)	,
(	3187	)	,
(	3184	)	,
(	3181	)	,
(	3178	)	,
(	3174	)	,
(	3171	)	,
(	3168	)	,
(	3165	)	,
(	3161	)	,
(	3158	)	,
(	3155	)	,
(	3152	)	,
(	3149	)	,
(	3145	)	,
(	3142	)	,
(	3139	)	,
(	3136	)	,
(	3133	)	,
(	3129	)	,
(	3126	)	,
(	3123	)	,
(	3120	)	,
(	3117	)	,
(	3114	)	,
(	3110	)	,
(	3107	)	,
(	3104	)	,
(	3101	)	,
(	3098	)	,
(	3095	)	,
(	3091	)	,
(	3088	)	,
(	3085	)	,
(	3082	)	,
(	3079	)	,
(	3076	)	,
(	3072	)	,
(	3069	)	,
(	3066	)	,
(	3063	)	,
(	3060	)	,
(	3057	)	,
(	3054	)	,
(	3050	)	,
(	3047	)	,
(	3044	)	,
(	3041	)	,
(	3038	)	,
(	3035	)	,
(	3032	)	,
(	3029	)	,
(	3026	)	,
(	3022	)	,
(	3019	)	,
(	3016	)	,
(	3013	)	,
(	3010	)	,
(	3007	)	,
(	3004	)	,
(	3001	)	,
(	2998	)	,
(	2995	)	,
(	2991	)	,
(	2988	)	,
(	2985	)	,
(	2982	)	,
(	2979	)	,
(	2976	)	,
(	2973	)	,
(	2970	)	,
(	2967	)	,
(	2964	)	,
(	2961	)	,
(	2958	)	,
(	2955	)	,
(	2951	)	,
(	2948	)	,
(	2945	)	,
(	2942	)	,
(	2939	)	,
(	2936	)	,
(	2933	)	,
(	2930	)	,
(	2927	)	,
(	2924	)	,
(	2921	)	,
(	2918	)	,
(	2915	)	,
(	2912	)	,
(	2909	)	,
(	2906	)	,
(	2903	)	,
(	2900	)	,
(	2897	)	,
(	2894	)	,
(	2891	)	,
(	2888	)	,
(	2885	)	,
(	2882	)	,
(	2879	)	,
(	2876	)	,
(	2873	)	,
(	2870	)	,
(	2867	)	,
(	2864	)	,
(	2861	)	,
(	2858	)	,
(	2855	)	,
(	2852	)	,
(	2849	)	,
(	2846	)	,
(	2843	)	,
(	2840	)	,
(	2837	)	,
(	2834	)	,
(	2831	)	,
(	2828	)	,
(	2825	)	,
(	2822	)	,
(	2819	)	,
(	2816	)	,
(	2813	)	,
(	2810	)	,
(	2807	)	,
(	2804	)	,
(	2802	)	,
(	2799	)	,
(	2796	)	,
(	2793	)	,
(	2790	)	,
(	2787	)	,
(	2784	)	,
(	2781	)	,
(	2778	)	,
(	2775	)	,
(	2772	)	,
(	2769	)	,
(	2766	)	,
(	2763	)	,
(	2761	)	,
(	2758	)	,
(	2755	)	,
(	2752	)	,
(	2749	)	,
(	2746	)	,
(	2743	)	,
(	2740	)	,
(	2737	)	,
(	2734	)	,
(	2732	)	,
(	2729	)	,
(	2726	)	,
(	2723	)	,
(	2720	)	,
(	2717	)	,
(	2714	)	,
(	2711	)	,
(	2708	)	,
(	2706	)	,
(	2703	)	,
(	2700	)	,
(	2697	)	,
(	2694	)	,
(	2691	)	,
(	2688	)	,
(	2686	)	,
(	2683	)	,
(	2680	)	,
(	2677	)	,
(	2674	)	,
(	2671	)	,
(	2668	)	,
(	2666	)	,
(	2663	)	,
(	2660	)	,
(	2657	)	,
(	2654	)	,
(	2651	)	,
(	2649	)	,
(	2646	)	,
(	2643	)	,
(	2640	)	,
(	2637	)	,
(	2635	)	,
(	2632	)	,
(	2629	)	,
(	2626	)	,
(	2623	)	,
(	2620	)	,
(	2618	)	,
(	2615	)	,
(	2612	)	,
(	2609	)	,
(	2607	)	,
(	2604	)	,
(	2601	)	,
(	2598	)	,
(	2595	)	,
(	2593	)	,
(	2590	)	,
(	2587	)	,
(	2584	)	,
(	2581	)	,
(	2579	)	,
(	2576	)	,
(	2573	)	,
(	2570	)	,
(	2568	)	,
(	2565	)	,
(	2562	)	,
(	2559	)	,
(	2557	)	,
(	2554	)	,
(	2551	)	,
(	2548	)	,
(	2546	)	,
(	2543	)	,
(	2540	)	,
(	2537	)	,
(	2535	)	,
(	2532	)	,
(	2529	)	,
(	2526	)	,
(	2524	)	,
(	2521	)	,
(	2518	)	,
(	2516	)	,
(	2513	)	,
(	2510	)	,
(	2507	)	,
(	2505	)	,
(	2502	)	,
(	2499	)	,
(	2497	)	,
(	2494	)	,
(	2491	)	,
(	2488	)	,
(	2486	)	,
(	2483	)	,
(	2480	)	,
(	2478	)	,
(	2475	)	,
(	2472	)	,
(	2470	)	,
(	2467	)	,
(	2464	)	,
(	2461	)	,
(	2459	)	,
(	2456	)	,
(	2453	)	,
(	2451	)	,
(	2448	)	,
(	2445	)	,
(	2443	)	,
(	2440	)	,
(	2437	)	,
(	2435	)	,
(	2432	)	,
(	2429	)	,
(	2427	)	,
(	2424	)	,
(	2422	)	,
(	2419	)	,
(	2416	)	,
(	2414	)	,
(	2411	)	,
(	2408	)	,
(	2406	)	,
(	2403	)	,
(	2400	)	,
(	2398	)	,
(	2395	)	,
(	2393	)	,
(	2390	)	,
(	2387	)	,
(	2385	)	,
(	2382	)	,
(	2379	)	,
(	2377	)	,
(	2374	)	,
(	2372	)	,
(	2369	)	,
(	2366	)	,
(	2364	)	,
(	2361	)	,
(	2359	)	,
(	2356	)	,
(	2353	)	,
(	2351	)	,
(	2348	)	,
(	2346	)	,
(	2343	)	,
(	2340	)	,
(	2338	)	,
(	2335	)	,
(	2333	)	,
(	2330	)	,
(	2328	)	,
(	2325	)	,
(	2322	)	,
(	2320	)	,
(	2317	)	,
(	2315	)	,
(	2312	)	,
(	2310	)	,
(	2307	)	,
(	2305	)	,
(	2302	)	,
(	2299	)	,
(	2297	)	,
(	2294	)	,
(	2292	)	,
(	2289	)	,
(	2287	)	,
(	2284	)	,
(	2282	)	,
(	2279	)	,
(	2277	)	,
(	2274	)	,
(	2272	)	,
(	2269	)	,
(	2266	)	,
(	2264	)	,
(	2261	)	,
(	2259	)	,
(	2256	)	,
(	2254	)	,
(	2251	)	,
(	2249	)	,
(	2246	)	,
(	2244	)	,
(	2241	)	,
(	2239	)	,
(	2236	)	,
(	2234	)	,
(	2231	)	,
(	2229	)	,
(	2226	)	,
(	2224	)	,
(	2221	)	,
(	2219	)	,
(	2216	)	,
(	2214	)	,
(	2211	)	,
(	2209	)	,
(	2207	)	,
(	2204	)	,
(	2202	)	,
(	2199	)	,
(	2197	)	,
(	2194	)	,
(	2192	)	,
(	2189	)	,
(	2187	)	,
(	2184	)	,
(	2182	)	,
(	2179	)	,
(	2177	)	,
(	2175	)	,
(	2172	)	,
(	2170	)	,
(	2167	)	,
(	2165	)	,
(	2162	)	,
(	2160	)	,
(	2157	)	,
(	2155	)	,
(	2153	)	,
(	2150	)	,
(	2148	)	,
(	2145	)	,
(	2143	)	,
(	2141	)	,
(	2138	)	,
(	2136	)	,
(	2133	)	,
(	2131	)	,
(	2128	)	,
(	2126	)	,
(	2124	)	,
(	2121	)	,
(	2119	)	,
(	2116	)	,
(	2114	)	,
(	2112	)	,
(	2109	)	,
(	2107	)	,
(	2104	)	,
(	2102	)	,
(	2100	)	,
(	2097	)	,
(	2095	)	,
(	2093	)	,
(	2090	)	,
(	2088	)	,
(	2085	)	,
(	2083	)	,
(	2081	)	,
(	2078	)	,
(	2076	)	,
(	2074	)	,
(	2071	)	,
(	2069	)	,
(	2066	)	,
(	2064	)	,
(	2062	)	,
(	2059	)	,
(	2057	)	,
(	2055	)	,
(	2052	)	,
(	2050	)	,
(	2048	)	,
(	2045	)	,
(	2043	)	,
(	2041	)	,
(	2038	)	,
(	2036	)	,
(	2034	)	,
(	2031	)	,
(	2029	)	,
(	2027	)	,
(	2024	)	,
(	2022	)	,
(	2020	)	,
(	2017	)	,
(	2015	)	,
(	2013	)	,
(	2011	)	,
(	2008	)	,
(	2006	)	,
(	2004	)	,
(	2001	)	,
(	1999	)	,
(	1997	)	,
(	1994	)	,
(	1992	)	,
(	1990	)	,
(	1988	)	,
(	1985	)	,
(	1983	)	,
(	1981	)	,
(	1978	)	,
(	1976	)	,
(	1974	)	,
(	1972	)	,
(	1969	)	,
(	1967	)	,
(	1965	)	,
(	1962	)	,
(	1960	)	,
(	1958	)	,
(	1956	)	,
(	1953	)	,
(	1951	)	,
(	1949	)	,
(	1947	)	,
(	1944	)	,
(	1942	)	,
(	1940	)	,
(	1938	)	,
(	1935	)	,
(	1933	)	,
(	1931	)	,
(	1929	)	,
(	1926	)	,
(	1924	)	,
(	1922	)	,
(	1920	)	,
(	1917	)	,
(	1915	)	,
(	1913	)	,
(	1911	)	,
(	1909	)	,
(	1906	)	,
(	1904	)	,
(	1902	)	,
(	1900	)	,
(	1897	)	,
(	1895	)	,
(	1893	)	,
(	1891	)	,
(	1889	)	,
(	1886	)	,
(	1884	)	,
(	1882	)	,
(	1880	)	,
(	1878	)	,
(	1875	)	,
(	1873	)	,
(	1871	)	,
(	1869	)	,
(	1867	)	,
(	1865	)	,
(	1862	)	,
(	1860	)	,
(	1858	)	,
(	1856	)	,
(	1854	)	,
(	1851	)	,
(	1849	)	,
(	1847	)	,
(	1845	)	,
(	1843	)	,
(	1841	)	,
(	1838	)	,
(	1836	)	,
(	1834	)	,
(	1832	)	,
(	1830	)	,
(	1828	)	,
(	1826	)	,
(	1823	)	,
(	1821	)	,
(	1819	)	,
(	1817	)	,
(	1815	)	,
(	1813	)	,
(	1811	)	,
(	1808	)	,
(	1806	)	,
(	1804	)	,
(	1802	)	,
(	1800	)	,
(	1798	)	,
(	1796	)	,
(	1793	)	,
(	1791	)	,
(	1789	)	,
(	1787	)	,
(	1785	)	,
(	1783	)	,
(	1781	)	,
(	1779	)	,
(	1777	)	,
(	1774	)	,
(	1772	)	,
(	1770	)	,
(	1768	)	,
(	1766	)	,
(	1764	)	,
(	1762	)	,
(	1760	)	,
(	1758	)	,
(	1756	)	,
(	1754	)	,
(	1751	)	,
(	1749	)	,
(	1747	)	,
(	1745	)	,
(	1743	)	,
(	1741	)	,
(	1739	)	,
(	1737	)	,
(	1735	)	,
(	1733	)	,
(	1731	)	,
(	1729	)	,
(	1727	)	,
(	1725	)	,
(	1722	)	,
(	1720	)	,
(	1718	)	,
(	1716	)	,
(	1714	)	,
(	1712	)	,
(	1710	)	,
(	1708	)	,
(	1706	)	,
(	1704	)	,
(	1702	)	,
(	1700	)	,
(	1698	)	,
(	1696	)	,
(	1694	)	,
(	1692	)	,
(	1690	)	,
(	1688	)	,
(	1686	)	,
(	1684	)	,
(	1682	)	,
(	1680	)	,
(	1678	)	,
(	1676	)	,
(	1674	)	,
(	1672	)	,
(	1670	)	,
(	1668	)	,
(	1666	)	,
(	1664	)	,
(	1662	)	,
(	1660	)	,
(	1658	)	,
(	1656	)	,
(	1654	)	,
(	1652	)	,
(	1650	)	,
(	1648	)	,
(	1646	)	,
(	1644	)	,
(	1642	)	,
(	1640	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1632	)	,
(	1630	)	,
(	1628	)	,
(	1626	)	,
(	1624	)	,
(	1622	)	,
(	1620	)	,
(	1618	)	,
(	1616	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1600	)	,
(	1598	)	,
(	1596	)	,
(	1594	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1583	)	,
(	1581	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1566	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1550	)	,
(	1548	)	,
(	1546	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1447	)	,
(	1445	)	,
(	1443	)	,
(	1441	)	,
(	1439	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1385	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1378	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1352	)	,
(	1350	)	,
(	1348	)	,
(	1347	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1321	)	,
(	1319	)	,
(	1318	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1311	)	,
(	1309	)	,
(	1308	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1281	)	,
(	1280	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1263	)	,
(	1262	)	,
(	1260	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1250	)	,
(	1249	)	,
(	1247	)	,
(	1246	)	,
(	1244	)	,
(	1242	)	,
(	1241	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1234	)	,
(	1233	)	,
(	1231	)	,
(	1230	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1190	)	,
(	1189	)	,
(	1187	)	,
(	1186	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1178	)	,
(	1176	)	,
(	1175	)	,
(	1173	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1166	)	,
(	1164	)	,
(	1163	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1155	)	,
(	1154	)	,
(	1152	)	,
(	1151	)	,
(	1149	)	,
(	1148	)	,
(	1146	)	,
(	1145	)	,
(	1143	)	,
(	1142	)	,
(	1140	)	,
(	1139	)	,
(	1137	)	,
(	1136	)	,
(	1134	)	,
(	1133	)	,
(	1131	)	,
(	1130	)	,
(	1128	)	,
(	1127	)	,
(	1125	)	,
(	1124	)	,
(	1122	)	,
(	1121	)	,
(	1119	)	,
(	1118	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1110	)	,
(	1109	)	,
(	1107	)	,
(	1106	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1100	)	,
(	1099	)	,
(	1097	)	,
(	1096	)	,
(	1094	)	,
(	1093	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1087	)	,
(	1086	)	,
(	1084	)	,
(	1083	)	,
(	1081	)	,
(	1080	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1074	)	,
(	1073	)	,
(	1071	)	,
(	1070	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1064	)	,
(	1063	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1057	)	,
(	1056	)	,
(	1054	)	,
(	1053	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1047	)	,
(	1046	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1036	)	,
(	1035	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1029	)	,
(	1028	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1018	)	,
(	1017	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	999	)	,
(	998	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	799	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	751	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	319	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	316	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	311	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	309	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	307	)	,
(	307	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	305	)	,
(	305	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	303	)	,
(	303	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	301	)	,
(	301	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	298	)	,
(	298	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	295	)	,
(	295	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	292	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	289	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	285	)	,
(	285	)	,
(	285	)	,
(	284	)	,
(	284	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	282	)	,
(	282	)	,
(	282	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	269	)	,
(	269	)	,
(	269	)	,
(	268	)	,
(	268	)	,
(	268	)	,
(	267	)	,
(	267	)	,
(	267	)	,
(	267	)	,
(	266	)	,
(	266	)	,
(	266	)	,
(	265	)	,
(	265	)	,
(	265	)	,
(	264	)	,
(	264	)	,
(	264	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	262	)	,
(	262	)	,
(	262	)	,
(	261	)	,
(	261	)	,
(	261	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	259	)	,
(	259	)	,
(	259	)	,
(	258	)	,
(	258	)	,
(	258	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	256	)	,
(	256	)	,
(	256	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	254	)	,
(	254	)	,
(	254	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	252	)	,
(	252	)	,
(	252	)	,
(	251	)	,
(	251	)	,
(	251	)	,
(	251	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	249	)	,
(	249	)	,
(	249	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	245	)	,
(	245	)	,
(	245	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	229	)	,
(	229	)	,
(	229	)	,
(	229	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	227	)	,
(	227	)	,
(	227	)	,
(	227	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	163	)	




);


end package LUT_pkg;
